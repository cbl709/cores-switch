`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:24:31 12/12/2012 
// Design Name: 
// Module Name:    pulse_detection 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "uart_defines.v"
module pulse_detection(
								clk,
								pwm,
								io
								);
input clk;
input pwm;
output io;	

parameter Period = `OSC;		// use 14.7456MHZ OSC,0.001s	


reg [31:0] time_counter     =32'h0000;
reg [31:0] rise_match_time  =32'h0000;
reg [31:0] fall_match_time  =32'h0000;
reg io                      =1'b1; //��ʼ״̬��Ϊ��⵽��������ֹAB��������ʱ���ֻ���//edit in 2013-3-5

//////////////////detect 1khz 50% duty pwm signal ///////
reg pwm_d1                  =1'b0;
reg pwm_d2                  =1'b0;
reg start                   =1'b0;
reg start_d1                =1'b0; // start���һ��clk��ʱ�����жϲ����Ƿ���ȷ
always@ (posedge clk)
begin
 pwm_d1 <= pwm;
 pwm_d2 <= pwm_d1;
 start_d1 <= start;
end

wire rise_edge;
wire fall_edge;

reg freq_right             =1'b1;
reg duty_right             =1'b1;

assign rise_edge = pwm_d1&(~pwm_d2);
assign fall_edge = ~pwm_d1&pwm_d2;

always@ (posedge clk )
begin
	
	if(~start&rise_edge) begin	//��⵽�����أ�ʱ�Ӽ�����time_counter��ʼ��ʱ
		start				 <= 1;
		
	end
	
	if(start&fall_edge) begin  //��⵽�½��أ���¼�½���ʱ��
		fall_match_time <= time_counter;
	end
	
	if(start&rise_edge) begin  //��⵽�����أ�ֹͣ������������¼������ʱ��
		rise_match_time <= time_counter;
		start			<= 0;
	end
	 			
end

always@(posedge clk )
begin
		if(start)
		time_counter <= time_counter+1;
		if(~start_d1)
		time_counter <= 16'b0;
end

always@(posedge clk )
begin
    if(~start_d1) begin     // start�źŽ������ӳ�һ��clk�����clk�����жϲ��� //edit in 2013-3-5
		if( (rise_match_time>=(Period-50)) && (rise_match_time <= (Period+50)) )// ������������??��50 ?�clk
			freq_right <= 1;  // frequency is 1khz, right
		else
			freq_right <= 0;
			
		if( (fall_match_time>=(Period/2-50)) && (fall_match_time <= (Period/2+50)) )	
			duty_right <=1;  // duty is 50%,righ
		else
			duty_right <=0;	
	end  // end of start_d1
	
end
wire io_tmp;
assign io_tmp= freq_right&duty_right;

//// io_tmp==1 for more than DETECTION_TIME period, io=1;
reg [31:0] io_high_counter =32'h00000000;
reg [31:0] io_low_counter  =32'h00000000;
always@(posedge clk )
begin
		if(io_tmp) begin
			io_high_counter <= io_high_counter+1;
			io_low_counter <= 0;
			end
		else begin
			io_high_counter <= 0;
			io_low_counter <= io_low_counter+1;
		 end
		if(io_high_counter >= `DETECTION_TIME*Period) begin
			io <=1;
			io_high_counter <= 0;
		end
		if(io_low_counter >=  `DETECTION_TIME*Period) begin
			io <=0;
			io_low_counter <= 0;
		end
			
end

endmodule
